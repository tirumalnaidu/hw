
package nvdla_coverage_pkg;

    import uvm_pkg::*;
`include "uvm_macros.svh"

`include "project.vh"
   
    import csb_pkg::*;
    import nvdla_ral_pkg::*;

    `include "bit_toggle_cg.sv"
    `include "nvdla_coverage_define.sv"
    `include "nvdla_coverage_base.sv"
    `include "nvdla_coverage_conv.sv"
    `include "nvdla_coverage_sdp.sv"
    `include "nvdla_coverage_pdp.sv"
    `include "nvdla_coverage_cdp.sv"
    `include "nvdla_coverage_bdma.sv"
    `include "nvdla_coverage_rubik.sv"
    `include "nvdla_coverage_top.sv"

endpackage
